** Profile: "SCHEMATIC2-pro_up_2"  [ c:\users\meisam\appdata\roaming\spb_data\project1_elec2-PSpiceFiles\SCHEMATIC2\pro_up_2.sim ] 

** Creating circuit file "pro_up_2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../project1_elec2-pspicefiles/project1_elec2.lib" 
* From [PSPICE NETLIST] section of C:\Users\Meisam\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.008 0 1u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC2.net" 


.END
