** Profile: "project-pro_simu1"  [ c:\users\meisam\appdata\roaming\spb_data\project1_elec2-pspicefiles\project\pro_simu1.sim ] 

** Creating circuit file "pro_simu1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../project1_elec2-pspicefiles/project1_elec2.lib" 
* From [PSPICE NETLIST] section of C:\Users\Meisam\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.012 0 3u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\project.net" 


.END
